// ---------------------------------------------------------------------
//    Module:     Testbench for 32-bit 32:1 Mux
//    Author:     Alex Schendel and Kevin Hoser
//    Contact:    schendel21@up.edu and hoser21@up.edu
//    Date:       3/27/2020
//
//    All rights reserved
// ---------------------------------------------------------------------

`timescale 1ns / 1ns

module test_mux32_32;

wire [31:0] z;
reg [31:0] i0, i1, i2, i3, i4, i5, i6, i7, 
             i8, i9, i10, i11, i12, i13, i14, i15,
             i16, i17, i18, i19, i20, i21, i22, i23, 
             i24, i25, i26, i27, i28, i29, i30, i31;
reg [4:0] s;

mux32_32 dut (z, i0, i1, i2, i3, i4, i5, i6, i7, 
                    i8, i9, i10, i11, i12, i13, i14, i15,
                    i16, i17, i18, i19, i20, i21, i22, i23, 
                    i24, i25, i26, i27, i28, i29, i30, i31, s);

  
initial	// Test stimulus
  begin
    i0 = 32'h00000000;
    i1 = 32'h00000001;
    i2 = 32'h00000002;
    i3 = 32'h00000003;
    i4 = 32'h00000004;
    i5 = 32'h00000005;
    i6 = 32'h00000006;
    i7 = 32'h00000007;
    i8 = 32'h00000008;
    i9 = 32'h00000009;
    i10 = 32'h0000000A;
    i11 = 32'h0000000B;
    i12 = 32'h0000000C;
    i13 = 32'h0000000D;
    i14 = 32'h0000000E;
    i15 = 32'h0000000F;
    i16 = 32'h00000010;
    i17 = 32'h00000011;
    i18 = 32'h00000012;
    i19 = 32'h00000013;
    i20 = 32'h00000014;
    i21 = 32'h00000015;
    i22 = 32'h00000016;
    i23 = 32'h00000017;
    i24 = 32'h00000018;
    i25 = 32'h00000019;
    i26 = 32'h0000001A;
    i27 = 32'h0000001B;
    i28 = 32'h0000001C;
    i29 = 32'h0000001D;
    i30 = 32'h0000001E;
    i31 = 32'h0000001F;
    s = 5'b00000;
    #10 s = 5'h01;
    #10 s = 5'h02;
    #10 s = 5'h03;
    #10 s = 5'h04;
    #10 s = 5'h05;
    #10 s = 5'h06;
    #10 s = 5'h07;
    #10 s = 5'h08;
    #10 s = 5'h09;
    #10 s = 5'h0A;
    #10 s = 5'h0B;
    #10 s = 5'h0C;
    #10 s = 5'h1E;
    #10 s = 5'h1F;
  end
    
endmodule  
